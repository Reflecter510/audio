BZh91AY&SY��� ���Ryg������?��� I  � @�P>�PNw+s@�2��F���4�b2d2��=CCF�JmG���F�4hA��� #@4S$"5=)�=L�Pѣ�  �   ��&�C##&��4@44�b $�"zL��0�d�MJ6�@4i��d�3H�CIV}�'BQI%Z@_�$�W�$H�	A�-]l�l�����EGiq
�����e�$E��(ʂ�eCl駃������"�]\�n�D�h��3��P����s��Ƒ����o����d��^����*�Pl���G�?-�Z�e�J��d������,��܌�o��/�e6.��IV�&�?n����EIay�`a�de���R#�;�^6�Z���G VH����X�5e`��g%]��4k�sk�h6`o4���bI��K�r'kَd�'�Il̥��N�UJ��0��XZI=Β$(BA���� �j�2��8��!*X8��#���D|F(�Ys�m`͂��[\��(T���E���C����؛�Ҝx��������LR�db���4G��U"A떛JVg>�yCz�nB8�&<(��y�s"�2e���@<#��A�8zB����&AQm!85ֈF��	6&��&O �1<d��Ť���.�o8Di��r)�F?K^&�,���cG
`�@1�*Ϋ��P�M5,��M¨�C�u�A0W�;�-d&��u��U�e	A@n�����
��|�̘=��pC\���nx�$L�(C�����;]�ɵeь�I*��r��ע��82�RKR+A�X.��ҭi&�������<�ɠ'�@6�rJjG��w,��/�)���i�c�D��uQ�6p�&1dGV,
,v�\�\;��.@,�K����ZA��o�*W�:bQ�PI�0Y�Ԁ@�':�l� ��!�ÿ*S��C�����U�}��.�DwSL�h���&G$2"&�g�!���#� ���6�NQ�.lg���ٖ�;J�fN"�I~��1hi�Hj0c+�b:�<%��%��w�+��Z]�F�#��:�2d��N���3I�T(��:,K�����P��C!�c�hs@ ڰ0jq �{r��@�R�6�*�)�&�}[B����"�",�b6�n��{؁�}O�@����`���avd2<_+����P�6�1�F,2�I��&�Ŗ�A�Qe!	z�T���w���xGlFaK�ü��i� �y�w���m���ܑN$><C� 